`timescale 1ns/1ps

module cpu (
    input clk, rst
);

endmodule